module johnson_counter();
  
endmodule