module hello_world;

initial
begin
  // This is a single line comment

  /*
  * This is 
  * a multi-line comment
  */

 $display("Hello World\n");
 $finish;
end

endmodule
